`timescale 1ns/1ps
// Wrapper to expose a dedicated Am95xx P2 scalar test target.
module tb_am95xx_p2_scalar;
  tb_am9513_scalar u_scalar();
endmodule
