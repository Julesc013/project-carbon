`timescale 1ns/1ps

module tb_z85_directed;
  tb_z85 #(.RUN_ZEX(1'b0)) u_tb();
endmodule
