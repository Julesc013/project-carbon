`timescale 1ns/1ps

module tb_z85_zex;
  tb_z85 #(.RUN_ZEX(1'b1)) u_tb();
endmodule
