`timescale 1ns/1ps

module tb_z90_directed;
  tb_z90 u_tb();
endmodule
