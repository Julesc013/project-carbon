`timescale 1ns/1ps
// Wrapper to expose a dedicated Am95xx P4 tensor test target.
module tb_am95xx_p4_tensor;
  tb_am9515_tensor u_tensor();
endmodule
