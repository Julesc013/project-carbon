`timescale 1ns/1ps
// Wrapper to expose a dedicated Am95xx P0 test target.
module tb_am95xx_p0;
  tb_am9513_scalar u_scalar();
endmodule
