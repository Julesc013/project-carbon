`timescale 1ns/1ps
// Wrapper to expose a dedicated Am95xx P3 vector test target.
module tb_am95xx_p3_vector;
  tb_am9514_vector u_vector();
endmodule
